library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity decoder is

	PORT(
		in_inst : std_logic_vector;
		out_inst : std_logic_vector
	);

end decoder;

architecture Behavioral of decoder is

begin

	


end Behavioral;

