library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity mux is

	PORT (
		data1 : std_logic_vector(15 downto 0);
		data2 : std_logic_vector(15 downto 0)
	);

end mux;

architecture Behavioral of mux is

begin

	process
	
		begin
		
			
		
	end process;


end Behavioral;

